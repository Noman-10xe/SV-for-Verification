/////////////////////////////////////////////////////////////////////
//   															   //
//   		  		   Scoreboard Class                            //
//                                                                 //
/////////////////////////////////////////////////////////////////////
//                                                                 //
//             Copyright (C) 2024 10xEngineers 	                   //
//             www.10xengineers.ai                                 //
//                                                                 //
/////////////////////////////////////////////////////////////////////
// FILE NAME      : scoreboard.sv
// AUTHOR         : Noman Rafiq
// AUTHOR'S EMAIL : noman.rafiq@10xengineers.ai
// ------------------------------------------------------------------
// RELEASE HISTORY													 
// ------------------------------------------------------------------
// VERSION DATE        	AUTHOR         								 
// 1.0     2024-Sep-27  Noman Rafiq 						 		 
// ------------------------------------------------------------------


// Include Function Definitions
`include "others.sv"

//////////////////////////////////////////////////////////////////
//
// Class Definition
//
class scoreboard;  
  
  //////////////////////////////////////////////////////////////////
  //
  // Declarations
  //
  mailbox mon2sco;		// Mailbox
  int no_transactions;	// To Track Number of Transactions
  bit	prev_reset;		// Stores Previous Value of Reset
  
  
  
  //////////////////////////////////////////////////////////////////
  //
  // Constructor
  //
  function new(mailbox mon2sco);
    this.mon2sco = mon2sco;
    $readmemh("memory_init.mem", mem);										// Initialize Memory to a Known State
    
    /*																
     *	Only Enable rd_mem.mem if you are trying to run rd_test.    
     *																
     *	"rd_mem.mem" is a memory initialized to randomly generated	
	 *	numbers so we can verify read operations.                  	
     *                                                             	
     *	[NOTE] :: Make sure to provide the DUT with the same 	  	
     *	Memory as Scoreboard for correct configuration. (INIT_FILE)	
     */

	//$readmemh("rd_mem.mem", mem);										// For rd_test Only
  
  endfunction
  
  
  //////////////////////////////////////////////////////////////////
  //
  // Main Method
  //
  
  // Stores HWDATA and compare HRDATA with the stored data
  task main();
  transaction t;
  forever begin
    mon2sco.get(t);

  	// Check if Reset is Asserted
    if (!t.HRESETn && prev_reset) begin
      $display("Local Memory Reset");
      $readmemh("memory_init.mem", mem);								// Initialize Memory to a Known State upon reset
    end else begin
      
      if (t.HREADY == 1'b1) begin 										// Check if Master is READY
        $display("[SCB] :: Transfer Can be Initiated");

        if (t.HPROT == 4'd1) begin 										// Checks if HPROT == 1
          $display("[SCB] :: Protection is set to DATA ACCESS Only");

          if (t.HSEL == 1'b1) begin 									// Check if Slave is Selected for Transfer
            $display("[SCB] :: Slave has been Selected");

            									
            if (t.HPROT == 4'd1) begin									// Perform Transfers when Data Access is Enabled
              
              
              //////////////////////////////////////////////////////////////////
              //
              // IDLE Transfer
              if (t.HTRANS == 2'b00) begin
                if (t.HRESP == 1'b0) 									// Checks for IDLE Transfer
                  $display("[SCB-PASS] :: IDLE TRANSFER :: SLAVE has provided with Zero Wait States (Okay Status).");
                else
                  $display("[SCB-FAIL] :: IDLE TRANSFER :: SLAVE has provided with Error Response.");
              end 

              
              //////////////////////////////////////////////////////////////////
              //
              // BUSY Transfer
              else if (t.HTRANS == 2'b01) begin
                if (t.HRESP == 1'b0) 									// Checks for BUSY Transfer
                  $display("[SCB-PASS] :: BUSY TRANSFER :: SLAVE has provided with Zero Wait States (Okay Status).");
                else
                  $display("[SCB-FAIL] :: BUSY TRANSFER :: SLAVE has provided with Error Response.");
              end 

              
              //////////////////////////////////////////////////////////////////
              //
              // NONSEQ Transfer
              else if (t.HTRANS == 2'b10) begin 						// Checks for NONSEQ Transfer
                if (t.HWRITE == 1'b1) WRITE(t); 						// NONSEQ Write
                else if (t.HWRITE == 1'b0) READ(t); 					// NONSEQ Read
              end 
              
			  
              //////////////////////////////////////////////////////////////////
              //
              // SEQ Transfer
              else if (t.HTRANS == 2'b11) begin 						// Checks for SEQ Transfer
                if (t.HWRITE == 1'b1) WRITE(t); 						// SEQ Write
                else if (t.HWRITE == 1'b0) READ(t); 					// SEQ Read
              end 
              
              else begin
                $display("[SCB-FAIL] :: HPROT should have been set to (1) => DATA ACCESS ONLY");
              end
            end

            
            //////////////////////////////////////////////////////////////////
  			//
  			// BURST CASE
  			//
            
//             if (t.HBURST == 3'd0 || t.HBURST == 3'd2 || t.HBURST == 3'd3) begin // Check the Type of BURST
//               																	// 0 (Single BURST), 2 (WRAP4), 3 (INCR4 BURST)
//               // SINGLE BURST
//               if (t.HBURST == 3'd0) begin
//                 if (t.HWRITE == 1) WRITE(t);
//                 else if (t.HWRITE == 0) READ(t);
//                 $display("[SCB] :: SINGLE BURST TRANSFER");
//               end 
              
//               // WRAP4 BURST
//               else if (t.HBURST == 3'd2) begin
//                 if (t.HWRITE == 1) WRITE(t);
//                 else if (t.HWRITE == 0) READ(t);
//                 $display("[SCB] :: 4-beat WRAPPING BURST");
//               end 
              
//               // INCR4 BURST
//               else if (t.HBURST == 3'd3) begin
//                 if (t.HWRITE == 1) WRITE(t);
//                 else if (t.HWRITE == 0) READ(t);
//                 $display("[SCB] :: 4-beat INCREMENTING BURST");
//               end
//             end
          end
        end
        no_transactions++;
      end 
        
        else begin
          
          // Check for Wait State
          if (t.HREADYOUT == 1'b0) begin
            $display("[SCB] :: Slave has inserted Wait States");
          end
          
          // Check if Slave is Connected
          if (t.HSEL == 1'b0) begin
            $display("[SCB] :: Slave has not been Connected");
          end
          
          no_transactions++;
        end 
      end
    
    prev_reset = t.HRESETn;
    
//     $display("--------- [Scoreboard - %0d] Debug Data  ------", no_transactions);
//     $display("\t HADDR 		= 0x%0h", t.HADDR);
//     $display("\t HWDATA 	= 0x%0h", t.HWDATA);
//     $display("\t HRDATA 	= 0x%0h", t.HRDATA);
//     $display("\t HWRITE		= %0b", t.HWRITE);
//     $display("\t HSIZE 		= %0b", t.HSIZE);
//     $display("\t HBURST 	= %0b", t.HBURST);
//     $display("\t HPROT 		= %0b", t.HPROT);
//     $display("\t HTRANS		= %0b", t.HTRANS);
//     $display("\t HREADYOUT	= %0b", t.HREADYOUT);
//     $display("\t HREADY 	= %0b", t.HREADY);
//     $display("\t HRESP 		= %0b", t.HRESP);
//     $display("\t HSEL 		= %0b", t.HSEL);
//     $display("\t HRESETn 	= %0b", t.HRESETn);
//     $display("\t prev_reset = %0b", prev_reset);
//     $display("\t no_transactions 	= %0d", no_transactions);
//     $display("---------------------------------------------\n");
    end
endtask
endclass
